library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000"
        ); 
begin

   dataout <= memory(to_integer(unsigned(address))); 

end Behavioral; 
